module TopModule (
  input clk,
  input load,
  input [255:0] data,
  output reg [255:0] q
);
    reg [255:0] next_q;

    always @(posedge clk) begin
        if (load)
            q <= data;
        else
            q <= next_q;
    end

    integer i, j;
    always @* begin
        next_q = q;
        for (i = 0; i < 16; i++) begin
            for (j = 0; j < 16; j++) begin
                // Calculate the indices of the neighbors, wrapping around the edges
                int left = (j == 0) ? 15 : j - 1;
                int right = (j == 15) ? 0 : j + 1;
                int up = (i == 0) ? 15 : i - 1;
                int down = (i == 15) ? 0 : i + 1;

                // Calculate the linear index for neighbors
                int idx_ul = up * 16 + left;
                int idx_u = up * 16 + j;
                int idx_ur = up * 16 + right;
                int idx_l = i * 16 + left;
                int idx_r = i * 16 + right;
                int idx_dl = down * 16 + left;
                int idx_d = down * 16 + j;
                int idx_dr = down * 16 + right;
                int idx = i * 16 + j;

                // Count the number of alive neighbors
                int count = q[idx_ul] + q[idx_u] + q[idx_ur] + q[idx_l] + q[idx_r] + q[idx_dl] + q[idx_d] + q[idx_dr];

                // Apply the rules of the game
                case (q[idx_ul] + q[idx_u] + q[idx_ur] + q[idx_l] + q[idx_r] + q[idx_dl] + q[idx_d] + q[idx_dr])
                    2: next_q[idx] = q[idx]; // Stay the same
                    3: next_q[idx] = 1'b1;   // Become alive
                    default: next_q[idx] = 1'b0; // Become dead or stay dead
                endcase
            end
        end
    end
endmodule

/*
Illegal Assignment
*/

/*
The testbench simulated, but had errors. Please fix the module. The output of iverilog is as follows:
VCD info: dumpfile wave.vcd opened for output.
Hint: The first test case is a blinker (initial state = 256'h7). First mismatch occurred at cycle 2.
Hint:
Hint: Cycle 2:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000010
Hint:   q[239:224]     0000000000000000      0000000000000000
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000000      0000000000000000
Hint:   q[ 31: 16]     0000000000000000      0000000000000010
Hint:   q[ 15:  0]     0000000000000110      0000000000000010
Hint:
Hint:

Hint: Cycle 3:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000000
Hint:   q[239:224]     0000000000000000      0000000000000000
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000000      0000000000000000
Hint:   q[ 31: 16]     0000000000000000      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000111
Hint:
Hint:

Hint: Cycle 4:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000010
Hint:   q[239:224]     0000000000000000      0000000000000000
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000000      0000000000000000
Hint:   q[ 31: 16]     0000000000000000      0000000000000010
Hint:   q[ 15:  0]     0000000000000110      0000000000000010
Hint:
Hint:

Hint: Cycle 5:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000000
Hint:   q[239:224]     0000000000000000      0000000000000000
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000000      0000000000000000
Hint:   q[ 31: 16]     0000000000000000      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000111
Hint:
Hint:

Hint: The second test case is a glider (initial state = 256'h000200010007). First mismatch occurred at cycle 2.
Hint:
Hint: Cycle 2:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000010
Hint:   q[239:224]     0000000000000000      0000000000000000
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000101
Hint:   q[ 15:  0]     0000000000000110      0000000000000011
Hint:
Hint:

Hint: Cycle 3:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000011
Hint:   q[239:224]     0000000000000000      0000000000000000
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000001
Hint:   q[ 15:  0]     0000000000000110      0000000000000101
Hint:
Hint:

Hint: Cycle 4:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000011
Hint:   q[239:224]     0000000000000000      0000000000000000
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000010
Hint:   q[ 15:  0]     0000000000000110      1000000000000001
Hint:
Hint:

Hint: Cycle 5:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      1000000000000011
Hint:   q[239:224]     0000000000000000      0000000000000000
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000001
Hint:   q[ 15:  0]     0000000000000110      1000000000000000
Hint:
Hint:

Hint: Cycle 6:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      1000000000000001
Hint:   q[239:224]     0000000000000000      0000000000000001
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      1000000000000010
Hint:
Hint:

Hint: Cycle 7:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      1000000000000010
Hint:   q[239:224]     0000000000000000      1000000000000001
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      1000000000000000
Hint:
Hint:

Hint: Cycle 8:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      1100000000000000
Hint:   q[239:224]     0000000000000000      1000000000000001
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000001
Hint:
Hint:

Hint: Cycle 9:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0100000000000000
Hint:   q[239:224]     0000000000000000      1100000000000001
Hint:   q[223:208]     0000000000000000      0000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      1000000000000000
Hint:
Hint:

Hint: Cycle 10:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0100000000000001
Hint:   q[239:224]     0000000000000000      1100000000000000
Hint:   q[223:208]     0000000000000000      1000000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000000
Hint:
Hint:

Hint: Cycle 11:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0100000000000000
Hint:   q[239:224]     0000000000000000      0100000000000001
Hint:   q[223:208]     0000000000000000      1100000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000000
Hint:
Hint:

Hint: Cycle 12:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      1000000000000000
Hint:   q[239:224]     0000000000000000      0110000000000000
Hint:   q[223:208]     0000000000000000      1100000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000000
Hint:
Hint:

Hint: Cycle 13:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0100000000000000
Hint:   q[239:224]     0000000000000000      0010000000000000
Hint:   q[223:208]     0000000000000000      1110000000000000
Hint:   q[207:192]     0000000000000000      0000000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000000
Hint:
Hint:

Hint: Cycle 14:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000000
Hint:   q[239:224]     0000000000000000      1010000000000000
Hint:   q[223:208]     0000000000000000      0110000000000000
Hint:   q[207:192]     0000000000000000      0100000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000000
Hint:
Hint:

Hint: Cycle 15:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000000
Hint:   q[239:224]     0000000000000000      0010000000000000
Hint:   q[223:208]     0000000000000000      1010000000000000
Hint:   q[207:192]     0000000000000000      0110000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000000
Hint:
Hint:

Hint: Cycle 16:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000000
Hint:   q[239:224]     0000000000000000      0100000000000000
Hint:   q[223:208]     0000000000000000      0011000000000000
Hint:   q[207:192]     0000000000000000      0110000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000000
Hint:
Hint:

Hint: Cycle 17:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000000
Hint:   q[239:224]     0000000000000000      0010000000000000
Hint:   q[223:208]     0000000000000000      0001000000000000
Hint:   q[207:192]     0000000000000000      0111000000000000
Hint:   q[191:176]     0000000000000000      0000000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000000
Hint:
Hint:

Hint: Cycle 18:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000000
Hint:   q[239:224]     0000000000000000      0000000000000000
Hint:   q[223:208]     0000000000000000      0101000000000000
Hint:   q[207:192]     0000000000000000      0011000000000000
Hint:   q[191:176]     0000000000000000      0010000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000000
Hint:
Hint:

Hint: Cycle 19:         Your game state       Reference game state
Hint:   q[255:240]     0000000000000000      0000000000000000
Hint:   q[239:224]     0000000000000000      0000000000000000
Hint:   q[223:208]     0000000000000000      0001000000000000
Hint:   q[207:192]     0000000000000000      0101000000000000
Hint:   q[191:176]     0000000000000000      0011000000000000
Hint:   q[175:160]     0000000000000000      0000000000000000
Hint:   q[159:144]     0000000000000000      0000000000000000
Hint:   q[143:128]     0000000000000000      0000000000000000
Hint:   q[127:112]     0000000000000000      0000000000000000
Hint:   q[111: 96]     0000000000000000      0000000000000000
Hint:   q[ 95: 80]     0000000000000000      0000000000000000
Hint:   q[ 79: 64]     0000000000000000      0000000000000000
Hint:   q[ 63: 48]     0000000000000000      0000000000000000
Hint:   q[ 47: 32]     0000000000000010      0000000000000000
Hint:   q[ 31: 16]     0000000000000001      0000000000000000
Hint:   q[ 15:  0]     0000000000000110      0000000000000000
Hint:
Hint:

./Execute_environment/testbench.sv:96: $finish called at 25116 (1ps)
Hint: Output 'q' has 5008 mismatches. First mismatch occurred at time 20.
Hint: Total mismatched samples is 5008 out of 5023 samples

Simulation finished at 25116 ps
Mismatches: 5008 in 5023 samples
*/