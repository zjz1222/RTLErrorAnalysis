
module TopModule (
  input [5:0] y,
  input w,
  output Y1,
  output Y3
);

assign Y1 = y[0] & ~y[1] | y[1] & ~y[2] | y[2] & ~y[4] | y[3] & ~w | y[4] & w;
assign Y3 = y[2] & ~y[3] | y[4] & w | y[5] & ~y[3];

endmodule
/*
Misinterpretation of Multimodal Data�� State Transition Diagram
*/
/*
The testbench simulated, but had errors. Please fix the module. The output of iverilog is as follows:
VCD info: dumpfile wave.vcd opened for output.
D:/MyVerilogDebugger/Dataset/dataset_verilog-eval-human/Prob091_2012_q2b_test.sv:45: $finish called at 3001 (1ps)
Hint: Output 'Y1' has 391 mismatches. First mismatch occurred at time 10.
Hint: Output 'Y3' has 253 mismatches. First mismatch occurred at time 10.
Hint: Total mismatched samples is 440 out of 600 samples

Simulation finished at 3001 ps
Mismatches: 440 in 600 samples

*/